interface mdio_if;
 logic tb_clk;
 logic clk;
 logic data;
 logic reset;
endinterface: mdio_if
