interface mdio_if;
 logic clk;
 logic data;
endinterface: mdio_if
