package mdio_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "mdio_driver.sv"
`include "mdio_env.sv"
`include "mdio_read_write_test.sv"

endpackage: mdio_pkg
