//kbilgund 
module top

endmodule 
