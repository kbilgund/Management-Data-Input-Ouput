interface mdio_if;
 logic tb_clk;
 logic clk;
 logic data;
endinterface: mdio_if
